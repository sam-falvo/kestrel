`default_nettype none
`timescale 1ns / 1ps
`include "asserts.vh"

module lsu_tb();
	reg	[11:0]	story_to;
	reg		fault_to;
	reg		clk_i, reset_i, we_i, nomem_i, hword_i, word_i;
	reg		dword_i;
	reg	[63:0]	addr_i, dat_i;
	reg	[1:0]	sel_i;

	wire		busy_o, rwe_o;
	wire	[63:0]	dat_o;

	wire	[63:0]	wbmadr_o;
	wire	[15:0]	wbmdat_o;
	wire		wbmwe_o, wbmstb_o;
	wire	[1:0]	wbmsel_o;
	reg		wbmack_i, wbmstall_i;
	reg	[15:0]	wbmdat_i;

	lsu ls(
		.clk_i(clk_i),
		.reset_i(reset_i),
		.addr_i(addr_i),
		.we_i(we_i),
		.nomem_i(nomem_i),
		.hword_i(hword_i),
		.word_i(word_i),
		.dword_i(dword_i),
		.busy_o(busy_o),
		.rwe_o(rwe_o),
		.dat_o(dat_o),
		.dat_i(dat_i),
		.sel_i(sel_i),

		.wbmadr_o(wbmadr_o),
		.wbmdat_o(wbmdat_o),
		.wbmwe_o(wbmwe_o),
		.wbmstb_o(wbmstb_o),
		.wbmsel_o(wbmsel_o),
		.wbmack_i(wbmack_i),
		.wbmstall_i(wbmstall_i),
		.wbmdat_i(wbmdat_i)
	);

	`STANDARD_FAULT
	`DEFASSERT0(busy, o)
	`DEFASSERT0(rwe, o)
	`DEFASSERT(dat, 63, o)
	`DEFASSERT(wbmadr, 63, o)
	`DEFASSERT(wbmdat, 15, o)
	`DEFASSERT(wbmsel, 1, o)
	`DEFASSERT0(wbmwe, o)
	`DEFASSERT0(wbmstb, o)

	always begin
		#5 clk_i <= ~clk_i;
	end

	task reset;
	begin
		reset_i <= 1;
		wait(~clk_i); wait(clk_i); #1;
		reset_i <= 0;
	end
	endtask

	initial begin
		$dumpfile("lsu.vcd");
		$dumpvars;

		{
		  wbmack_i, addr_i, dat_i, we_i, nomem_i, hword_i, word_i,
		  dword_i, clk_i, reset_i, story_to, fault_to, sel_i,
		  wbmstall_i
		} <= 0;

		wait(~clk_i); wait(clk_i); #1;

		reset;
		assert_busy(0);

		// Given that we're not accessing memory,
		// the LSU must pass the address through to the
		// register writeback stage.
		//
		// Note that we pass the address, and not the input
		// data, since that's the value generated by the CPU's
		// ALU (instruction execute) stage.

		story_to <= 12'h010;

		addr_i <= 64'h1122334455667788;
		dat_i <= 64'h7766554433221100;
		we_i <= 0;
		nomem_i <= 1;
		wait(~clk_i); wait(clk_i); #1;
		assert_dat(64'h1122334455667788);
		assert_rwe(1);

		story_to <= 12'h018;

		addr_i <= 64'h1122334455667788;
		dat_i <= 64'h7766554433221100;
		we_i <= 1;
		nomem_i <= 1;
		wait(~clk_i); wait(clk_i); #1;
		assert_dat(64'h1122334455667788);
		assert_rwe(1);

		we_i <= 0;

		// When idle, the LSU must disable writebacks to the register
		// file.

		story_to <= 12'h020;

		nomem_i <= 0;
		wait(~clk_i); wait(clk_i); #1;
		assert_rwe(0);

		// When writing a half-word to memory,
		// the LSU must initiate and wait for the complete
		// Wishbone transaction to complete.  Further, it must
		// disable register write-back.
		//
		// Note that the LSU performs both a read AND a write,
		// irrespective of the we_i signal.  It's up to the
		// external peripheral to respect the we_i signal.
		// Similarly, while the LSU "reads" data even during a
		// write transaction, the register writeback stage is
		// responsible for ignoring this value, as rd_i will be
		// forced to 0.

		story_to <= 12'h040;

		hword_i <= 1;
		addr_i <= 64'h1122334455667788;
		dat_i <= 64'h7766554433221100;
		we_i <= 1;
		wbmdat_i <= 16'hDEAD;
		sel_i <= 2'b11;

		wait(~clk_i); wait(clk_i); #1;

		hword_i <= 0;
		we_i <= 0;

		assert_busy(1);
		assert_wbmadr(64'h1122334455667788);
		assert_wbmdat(16'h1100);
		assert_wbmwe(1);
		assert_wbmstb(1);
		assert_wbmsel(2'b11);
		assert_rwe(0);

		wait(~clk_i); wait(clk_i); #1;

		assert_busy(1);
		assert_wbmstb(0);
		assert_wbmsel(2'b00);
		assert_rwe(0);
		
		wbmack_i <= 1;

		wait(~clk_i); wait(clk_i); #1;

		assert_rwe(1);
		assert_dat(64'h000000000000DEAD);

		wbmack_i <= 0;

		// When writing a full-word to memory,
		// the LSU must initiate and wait for the complete
		// Wishbone transaction to complete.  In this case,
		// the transfer consists of two cycles (one for lowest
		// 16-bits, one for highest 16-bits).

		story_to <= 12'h050;

		word_i <= 1;
		addr_i <= 64'h1122334455667788;
		dat_i <= 64'h7766554433221100;
		we_i <= 1;
		wbmdat_i <= 16'hDEAD;

		wait(~clk_i); wait(clk_i); #1;

		word_i <= 0;
		we_i <= 0;

		assert_busy(1);
		assert_wbmadr(64'h112233445566778A);
		assert_wbmdat(16'h3322);
		assert_wbmwe(1);
		assert_wbmstb(1);
		assert_wbmsel(2'b11);
		assert_rwe(0);

		wait(~clk_i); wait(clk_i); #1;

		assert_busy(1);
		assert_wbmadr(64'h1122334455667788);
		assert_wbmdat(16'h1100);
		assert_wbmwe(1);
		assert_wbmstb(1);
		assert_wbmsel(2'b11);
		assert_rwe(0);

		wait(~clk_i); wait(clk_i); #1;

		assert_busy(1);
		assert_wbmstb(0);
		assert_wbmsel(2'b00);
		assert_rwe(0);
		
		wbmack_i <= 1;
		wbmdat_i <= 16'hDEAD;

		wait(~clk_i); wait(clk_i); #1;

		wbmdat_i <= 16'hBEEF;

		wait(~clk_i); wait(clk_i); #1;

		assert_rwe(1);
		assert_dat(64'h00000000DEADBEEF);

		wbmack_i <= 0;

		// When writing a double-word to memory,
		// the LSU must initiate and wait for the complete
		// Wishbone transaction to complete.  In this case,
		// the transfer consists of four cycles.

		story_to <= 12'h060;

		dword_i <= 1;
		addr_i <= 64'h1122334455667788;
		dat_i <= 64'h7766554433221100;
		we_i <= 1;

		wait(~clk_i); wait(clk_i); #1;

		dword_i <= 0;
		we_i <= 0;

		assert_busy(1);
		assert_wbmadr(64'h112233445566778E);
		assert_wbmdat(16'h7766);
		assert_wbmwe(1);
		assert_wbmstb(1);
		assert_wbmsel(2'b11);
		assert_rwe(0);

		wait(~clk_i); wait(clk_i); #1;

		assert_busy(1);
		assert_wbmadr(64'h112233445566778C);
		assert_wbmdat(16'h5544);
		assert_wbmwe(1);
		assert_wbmstb(1);
		assert_wbmsel(2'b11);
		assert_rwe(0);

		wait(~clk_i); wait(clk_i); #1;

		assert_busy(1);
		assert_wbmadr(64'h112233445566778A);
		assert_wbmdat(16'h3322);
		assert_wbmwe(1);
		assert_wbmstb(1);
		assert_wbmsel(2'b11);
		assert_rwe(0);

		wait(~clk_i); wait(clk_i); #1;

		assert_busy(1);
		assert_wbmadr(64'h1122334455667788);
		assert_wbmdat(16'h1100);
		assert_wbmwe(1);
		assert_wbmstb(1);
		assert_wbmsel(2'b11);
		assert_rwe(0);

		wait(~clk_i); wait(clk_i); #1;

		assert_busy(1);
		assert_wbmstb(0);
		assert_wbmsel(2'b00);
		assert_rwe(0);
		
		wbmack_i <= 1;
		wbmdat_i <= 16'hDEAD;

		wait(~clk_i); wait(clk_i); #1;

		wbmdat_i <= 16'hBEEF;

		wait(~clk_i); wait(clk_i); #1;

		wbmdat_i <= 16'h0BAD;

		wait(~clk_i); wait(clk_i); #1;

		wbmdat_i <= 16'hC0DE;

		wait(~clk_i); wait(clk_i); #1;

		assert_rwe(1);
		assert_dat(64'hDEADBEEF0BADC0DE);

		wbmack_i <= 0;

		// When writing individual bytes to memory,
		// yeah, you know the drill.  But this time, things
		// are a little different.
		//
		// Since half-words are the smallest unit of transfer
		// on any given clock cycle, the instruction decoder
		// must assert hword_i to commence the transfer (since a
		// single byte occupies only a single cycle).
		// However, sel_i must be either 2'b01 or 2'b10 to select
		// the appropriate byte lane.
		//
		// Also, in this condition, dat_i[7:0] is the source of
		// data to store (assuming we_i is set), while dat_o[7:0]
		// is always the data read back (if any), REGARDLESS of
		// which byte lane is enabled.

		// These tests exercise the lower byte.

		story_to <= 12'h080;

		hword_i <= 1;
		sel_i <= 2'b01;
		addr_i <= 64'h1122334455667788;
		dat_i <= 64'h77665544332211A5;
		we_i <= 1;
		wbmdat_i <= 16'hDEAD;

		wait(~clk_i); wait(clk_i); #1;

		hword_i <= 0;
		we_i <= 0;

		assert_busy(1);
		assert_wbmadr(64'h1122334455667788);
		assert_wbmdat(16'hA5A5);
		assert_wbmwe(1);
		assert_wbmstb(1);
		assert_wbmsel(2'b01);
		assert_rwe(0);

		wait(~clk_i); wait(clk_i); #1;

		assert_busy(1);
		assert_wbmstb(0);
		assert_wbmsel(2'b00);
		assert_rwe(0);
		
		wbmack_i <= 1;

		wait(~clk_i); wait(clk_i); #1;

		assert_rwe(1);
		assert_dat(64'h00000000000000AD);

		wbmack_i <= 0;

		// These tests exercise the upper byte.

		story_to <= 12'h088;

		hword_i <= 1;
		sel_i <= 2'b10;
		addr_i <= 64'h1122334455667788;
		dat_i <= 64'h77665544332211A5;
		we_i <= 1;
		wbmdat_i <= 16'hDEAD;

		wait(~clk_i); wait(clk_i); #1;

		hword_i <= 0;
		we_i <= 0;

		assert_busy(1);
		assert_wbmadr(64'h1122334455667788);
		assert_wbmdat(16'hA5A5);
		assert_wbmwe(1);
		assert_wbmstb(1);
		assert_wbmsel(2'b10);
		assert_rwe(0);

		wait(~clk_i); wait(clk_i); #1;

		assert_busy(1);
		assert_wbmstb(0);
		assert_wbmsel(2'b00);
		assert_rwe(0);
		
		wbmack_i <= 1;

		wait(~clk_i); wait(clk_i); #1;

		assert_rwe(1);
		assert_dat(64'h00000000000000DE);

		wbmack_i <= 0;

		// So far, all tests have exercised separated cycles for
		// bus commands and bus responses.  But, these operate over
		// independent sub-buses, so it should be possible to overlap
		// their operation.  The perfect, most ideal case would be
		// single-cycle response times.

		story_to <= 12'h0A0;

		dword_i <= 1;
		addr_i <= 64'h1122334455667788;
		dat_i <= 64'h7766554433221100;
		we_i <= 1;
		sel_i <= 2'b11;

		wait(~clk_i); wait(clk_i); #1;

		dword_i <= 0;
		we_i <= 0;

		assert_busy(1);
		assert_wbmadr(64'h112233445566778E);
		assert_wbmdat(16'h7766);
		assert_wbmwe(1);
		assert_wbmstb(1);
		assert_wbmsel(2'b11);
		assert_rwe(0);

		wbmack_i <= 1;
		wbmdat_i <= 16'hDEAD;

		wait(~clk_i); wait(clk_i); #1;

		assert_busy(1);
		assert_wbmadr(64'h112233445566778C);
		assert_wbmdat(16'h5544);
		assert_wbmwe(1);
		assert_wbmstb(1);
		assert_wbmsel(2'b11);
		assert_rwe(0);

		wbmdat_i <= 16'hBEEF;

		wait(~clk_i); wait(clk_i); #1;

		assert_busy(1);
		assert_wbmadr(64'h112233445566778A);
		assert_wbmdat(16'h3322);
		assert_wbmwe(1);
		assert_wbmstb(1);
		assert_wbmsel(2'b11);
		assert_rwe(0);

		wbmdat_i <= 16'hFEED;

		wait(~clk_i); wait(clk_i); #1;

		assert_busy(1);
		assert_wbmadr(64'h1122334455667788);
		assert_wbmdat(16'h1100);
		assert_wbmwe(1);
		assert_wbmstb(1);
		assert_wbmsel(2'b11);
		assert_rwe(0);

		wbmdat_i <= 16'hFACE;

		wait(~clk_i); wait(clk_i); #1;

		wbmack_i <= 0;

		assert_rwe(1);
		assert_dat(64'hDEADBEEFFEEDFACE);

		// The STALL_I signal is required to slow down the command-
		// phase of bus transactions.  We repeat a 64-bit transaction
		// here, but stall for 3 cycles mid-way.

		story_to <= 12'h0B0;

		dword_i <= 1;
		addr_i <= 64'h1122334455667788;
		dat_i <= 64'h7766554433221100;
		we_i <= 1;
		sel_i <= 2'b11;

		wait(~clk_i); wait(clk_i); #1;

		dword_i <= 0;
		we_i <= 0;

		assert_busy(1);
		assert_wbmadr(64'h112233445566778E);
		assert_wbmdat(16'h7766);
		assert_wbmwe(1);
		assert_wbmstb(1);
		assert_wbmsel(2'b11);
		assert_rwe(0);

		wait(~clk_i); wait(clk_i); #1;

		assert_busy(1);
		assert_wbmadr(64'h112233445566778C);
		assert_wbmdat(16'h5544);
		assert_wbmwe(1);
		assert_wbmstb(1);
		assert_wbmsel(2'b11);
		assert_rwe(0);

		wbmack_i <= 1;
		wbmdat_i <= 16'hFEED;

		wait(~clk_i); wait(clk_i); #1;

		assert_busy(1);
		assert_wbmadr(64'h112233445566778A);
		assert_wbmdat(16'h3322);
		assert_wbmwe(1);
		assert_wbmstb(1);
		assert_wbmsel(2'b11);
		assert_rwe(0);

		wbmstall_i <= 1;
		wbmack_i <= 0;

		wait(~clk_i); wait(clk_i); #1;

		assert_busy(1);
		assert_wbmadr(64'h112233445566778A);
		assert_wbmdat(16'h3322);
		assert_wbmwe(1);
		assert_wbmstb(1);
		assert_wbmsel(2'b11);
		assert_rwe(0);

		wbmstall_i <= 1;
		wbmack_i <= 0;

		wait(~clk_i); wait(clk_i); #1;

		assert_busy(1);
		assert_wbmadr(64'h112233445566778A);
		assert_wbmdat(16'h3322);
		assert_wbmwe(1);
		assert_wbmstb(1);
		assert_wbmsel(2'b11);
		assert_rwe(0);

		wbmstall_i <= 1;
		wbmack_i <= 0;

		wait(~clk_i); wait(clk_i); #1;

		assert_busy(1);
		assert_wbmadr(64'h112233445566778A);
		assert_wbmdat(16'h3322);
		assert_wbmwe(1);
		assert_wbmstb(1);
		assert_wbmsel(2'b11);
		assert_rwe(0);

		wbmstall_i <= 0;
		wbmack_i <= 1;
		wbmdat_i <= 16'hFACE;

		wait(~clk_i); wait(clk_i); #1;

		assert_busy(1);
		assert_wbmadr(64'h1122334455667788);
		assert_wbmdat(16'h1100);
		assert_wbmwe(1);
		assert_wbmstb(1);
		assert_wbmsel(2'b11);
		assert_rwe(0);

		wbmdat_i <= 16'h00C0;

		wait(~clk_i); wait(clk_i); #1;

		wbmdat_i <= 16'hFFEE;

		wait(~clk_i); wait(clk_i); #1;

		wbmack_i <= 0;
		wbmdat_i <= 0;

		assert_rwe(1);
		assert_dat(64'hFEEDFACE00C0FFEE);

		#100;
		$stop;
	end
endmodule

